top_cae.sv