CAE_srcs/parameters.sv